module fft_16_b4(
    input reg clk,
    input reg rst_n,
    input reg [17:0] x [15:0],
    output reg [17:0] Y [15:0]
);




endmodule