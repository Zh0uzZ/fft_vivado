module exp_resize #(
    parameter expWidth = 4
) (
    input [expWidth*32-1:0] input_exp,
    input [expWidth-1:0] max_exp,
    output [expWidth*32-1:0] output_exp
);
    

endmodule
